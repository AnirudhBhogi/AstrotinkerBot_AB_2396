
// reg_file.v - register file for single-cycle RISC-V CPU
//              (with 32 registers, each of 32 bits)
//              having two read ports, one write port
//              write port is synchronous, read ports are combinational
//              register 0 is hardwired to 0

module reg_file #(parameter DATA_WIDTH = 32) (
    input       clk,reset,
    input       wr_en,
    input       [4:0] rd_addr1, rd_addr2, wr_addr,
    input       [DATA_WIDTH-1:0] wr_data,
    output      [DATA_WIDTH-1:0] rd_data1, rd_data2,
	 output      flagr13_14
);

reg [DATA_WIDTH-1:0] reg_file_arr [0:31];
reg flag = 1'b0;
initial begin
	flag = 1'b0;
end
integer i;
initial begin
    for (i = 0; i < 32; i = i + 1) begin
        reg_file_arr[i] = 0;
    end
end

// register file write logic (synchronous)
always @(posedge clk) begin
//	if(!reset) begin
	if((^reset === 1'b0) && flag) begin
    if (wr_en) reg_file_arr[wr_addr] <= wr_data;
	 end
	else if((^reset===1'bz) || (^reset===1'b1) || (^reset===1'bx))
	begin flag <= 1'b1; end
end

// register file read logic (combinational)
assign rd_data1 = ( rd_addr1 != 0 ) ? reg_file_arr[rd_addr1] : 0;
assign rd_data2 = ( rd_addr2 != 0 ) ? reg_file_arr[rd_addr2] : 0;
assign flagr13_14 = (wr_addr==13 || wr_addr==14) ? 1 : 0;
endmodule
